* A Chain of 100 2-input AND Gates 
* Apply a pulse input to the chain and measure all timings
* Use the most recently characterized AND2 sub-circuit as the chain's
* basic element

* Either the normal version AND2 or the weak pin-B version AND2 included
.include ./working_and2_sckt.spice

* Configure the circuit and input signal settings
.param in_slope=0.04NS
.param last_stage_load_cap=0fF
.param every_10gates_cap=0fF

* Include the 100 stages chain circuit
.include ./and2_chain_sckt.spice

VCC vcc 0 1.1V
VIN vin 0 0 PULSE(1.1 0 0 {in_slope} {in_slope} 20NS 40NS)
* add source internal resistance to imitate real source
Rin vin drvin 10

* an inverter as the input driver
M1 vcc drvin 1 vcc p1 W=0.63u L=0.05u M=5
M2 1 drvin 0 0 n1 W=0.42u L=0.05u M=5
* a capacitor as the driver's fanout
Cdrvout 1 0 1fF

* two chains connected to the same node 1
X1 1 vcc 2 vcc AND2C100A
X2 vcc 1 3 vcc AND2C100B

C1 2 0 {last_stage_load_cap}
C2 3 0 {last_stage_load_cap}

.tran 0.01ns 50ns
.save V(1) V(2) V(3)

* if need all signals to debug
.save all

.measure tran tr_in TRIG V(1) VAL=0.33 RISE=2 TARG V(1) VAL=0.77 RISE=2
.measure tran tf_in TRIG V(1) VAL=0.77 FALL=1 TARG V(1) VAL=0.33 FALL=1
.measure tran tr_out_Ain TRIG V(2) VAL=0.33 RISE=2 TARG V(2) VAL=0.77 RISE=2
.measure tran tr_out_Bin TRIG V(3) VAL=0.33 RISE=2 TARG V(3) VAL=0.77 RISE=2
.measure tran tf_out_Ain TRIG V(2) VAL=0.77 FALL=1 TARG V(2) VAL=0.33 FALL=1
.measure tran tf_out_Bin TRIG V(3) VAL=0.77 FALL=1 TARG V(3) VAL=0.33 FALL=1
.measure tran tpdr_Ain TRIG V(1) VAL=0.55 RISE=2 TARG V(2) VAL=0.55 RISE=2
.measure tran tpdr_Bin TRIG V(1) VAL=0.55 RISE=2 TARG V(3) VAL=0.55 RISE=2
.measure tran tpdf_Ain TRIG V(1) VAL=0.55 FALL=1 TARG V(2) VAL=0.55 FALL=1
.measure tran tpdf_Bin TRIG V(1) VAL=0.55 FALL=1 TARG V(3) VAL=0.55 FALL=1

.end
