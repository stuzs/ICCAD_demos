* circuit of linear components plus diodes
dx 1 6 diode
dy 0 6 diode
rx 1 2 1
ry 2 3 1
rz 3 1 0.5
rg 1 0 1
ix 0 1 1
iz 0 3 1
r1 101 102 100
r2 102 0 10000
v1 101 0 5
d1 102 103 diode
d2 103 gnd diode
