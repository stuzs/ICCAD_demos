2-input AND Gate Cell Characterization Demo

.SUBCKT AND2 in1 in2 out VDD
* NODES: INPUT, INPUT, OUTPUT, VCC
* stage 1: PMOS VCC->M1//M2; NMOS M3--M4->GND
*  in1(pin A) controls M1 and M3
*  in2(pin B) controls M2 and M4
* stage 2: PMOS M5; NMOS M6
M1 net1 in1 Vdd Vdd p1 W=0.315u L=0.05u
M2 net1 in2 Vdd Vdd p1 W=0.315u L=0.05u
M3 net1 in1 net2 0 n1 W=0.21u L=0.05u
M4 0 in2 net2 0 n1 W=0.21u L=0.05u
M5 Vdd net1 out Vdd p1 W=0.63u L=0.05u
M6 out net1 0 0 n1 W=0.21u L=0.05u
.ENDS AND2

* use BSIM4 model with default parameter values,
* as if in a .lib TT library setting, and 
* ignore setting other FF, SS, FS, SF corners
.model n1 nmos level=54 version=4.8.0
.model p1 pmos level=54 version=4.8.0

* define the 2D-LUT index values,
* try changing parameter values in batch runs
.param slope=0.2NS
.param cap=10ff

VCC 4 0 DC 1.1V
VIN 1 0 DC 0 PULSE(0 1.1 0 {slope} {slope} 20NS 40NS)

* measure and compare V(1) and V(2) for timing characterization
X0 1 4 2 4 AND2
* but to characterize another input pin(i.e., switch A/B) we use
*X0 4 1 2 4 AND2

* the output load capacitor
CL 2 0 {cap}

.tran 0.001ns 100ns
.save V(1) V(2)
*.plot V(1) V(2)

* define level 30%->70% propagation delay
* and I choose the second rising edge to measure
.measure tran tr_in TRIG V(1) VAL=0.33 RISE=2 TARG V(1) VAL=0.77 RISE=2
.measure tran tr_out TRIG V(2) VAL=0.33 RISE=2 TARG V(2) VAL=0.77 RISE=2
.measure tran tdiff TRIG V(1) VAL=0.55 RISE=2 TARG V(2) VAL=0.55 RISE=2

*.control
*run
*.endc

.end
