* low pass filter
r1 1 2 10
r2 2 3 10
r3 3 0 10
z1 2 0 -100j
#z1 2 0 -10j
#z1 2 0 -1j
#z1 2 0 -0.1j
#z1 2 0 -0.01j
#z1 2 0 -0.001j
i1 0 1 1
