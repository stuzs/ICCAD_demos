* Example circuit shows LU decomposition on lecture slides
rx 1 2 1
ry 2 3 1
rz 3 1 0.5
rg 1 0 1
ix 0 1 1
iz 0 3 1
