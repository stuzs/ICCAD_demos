* 2-input AND Gate (AND2) Cell Characterization Demo
* Use alter method for batch running to generate NLDM 2-D timing table.

* Add an invert as driver to imitate real input driving condition.
* Add dirver loading capacitance to imitate driver's fan-out.
* Since the driving inverter will sharpen any slow input waveform, the
* driver's load capacitance is used to control the slew rate on test signal.

.include ./working_and2_sckt.spice

* define 3 parameters to control input waveform shape
* define another 1 parameter for output load
* all parameters changed during alterparam procedure
.param vin_slope=0.01NS
.param drv_load_cap=30fF
.param drv_M=10
.param out_load_cap=100fF

* input pulse voltage source with 10-Ohms internal resistance
VCC vcc 0 1.1V
VIN vin 0 0 PULSE(1.1 0 0 {vin_slope} {vin_slope} 20NS 40NS)
Rin vin drvin 10

* an inverter as the input driver, {drv_M} defines the multiplicity factor
M1 vcc drvin 1 vcc p1 W=0.63u L=0.05u M={drv_M}
M2 1 drvin 0 0 n1 W=0.42u L=0.05u M={drv_M}
* a capacitor as the driver's fanout
Cdrvout 1 0 {drv_load_cap}

*X1 for testing PIN A; node 1: input; node 2: output
X1 1 vcc 2 vcc AND2
CL1 2 0 {out_load_cap}

*X2 for testing PIN B; node 1: input; node 3: output
X2 vcc 1 3 vcc AND2
CL2 3 0 {out_load_cap}

*.tran 0.001n 100n
*.save all

* Use combinations of 3 input parameter values below.
* The purpose is to imitate input waveforms in more realistic
* working environment.
* For parameters vin_slope, drv_load_cap, drv_M
* 0.001n, 0.1f, 10 => fastest test signal, input slew: ~3ps
* 0.02n, 10f, 5 => input slew: ~7.5ps
* 0.05n, 20f, 3 => input slew: ~17.5ps
* 0.1n, 50f, 2 => input slew: ~41ps

* Output loading capacitances are chosen as below
* 0.3f, 2f, 10f, 50f

.control
compose input_param0 values 0.001n 0.02n 0.05n 0.3n
compose input_param1 values 0.1f 10f 20f 50f
compose input_param2 values 10 5 3 2
compose output_param values 0.3f 3f 20f 100f

foreach input_cond 0 1 2 3 
  foreach output_cond 0 1 2 3
    let pv1 = input_param0[$input_cond]
    let pv2 = input_param1[$input_cond]
    let pv3 = input_param2[$input_cond]
    let pv4 = output_param[$output_cond]
    set p1 = $&pv1
    set p2 = $&pv2
    set p3 = $&pv3
    set p4 = $&pv4
    echo ****************
    echo "AND2 cell characterization simulation with"
    echo "input condition case = $input_cond"
    echo "output condition case = $output_cond" 
    echo ****************
    alterparam vin_slope = $p1
    alterparam drv_load_cap = $p2
    alterparam drv_M = $p3
    alterparam out_load_cap = $p4
    reset $ reset is needed after alterparam
    tran 0.001ns 100ns
    run
*   define level 30%->70% propagation delay
*   and I choose the second rising edge and first falling edge to measure
    meas tran tr_in TRIG V(1) VAL=0.33 RISE=2 TARG V(1) VAL=0.77 RISE=2
    meas tran tf_in TRIG V(1) VAL=0.77 FALL=1 TARG V(1) VAL=0.33 FALL=1
    echo "out_load_cap        =  $p4"
    meas tran tr_out_Ain TRIG V(2) VAL=0.33 RISE=2 TARG V(2) VAL=0.77 RISE=2
    meas tran tr_out_Bin TRIG V(3) VAL=0.33 RISE=2 TARG V(3) VAL=0.77 RISE=2
    meas tran tf_out_Ain TRIG V(2) VAL=0.77 FALL=1 TARG V(2) VAL=0.33 FALL=1
    meas tran tf_out_Bin TRIG V(3) VAL=0.77 FALL=1 TARG V(3) VAL=0.33 FALL=1
    meas tran tpdr_Ain TRIG V(1) VAL=0.55 RISE=2 TARG V(2) VAL=0.55 RISE=2
    meas tran tpdr_Bin TRIG V(1) VAL=0.55 RISE=2 TARG V(3) VAL=0.55 RISE=2
    meas tran tpdf_Ain TRIG V(1) VAL=0.55 FALL=1 TARG V(2) VAL=0.55 FALL=1
    meas tran tpdf_Bin TRIG V(1) VAL=0.55 FALL=1 TARG V(3) VAL=0.55 FALL=1
  end
end
exit
.endc

.end
